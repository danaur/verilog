
module useaoi();
	wire a, b, c, d, f;

	AIO instance (a, b, c, d, f);
endmodule

